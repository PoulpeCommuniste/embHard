-- model.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity model is
	port (
		clk_clk                                : in    std_logic                     := '0';             --                             clk.clk
		lcd_dma_ctrl_0_conduit_end_lcd_d_c_n   : out   std_logic;                                        --      lcd_dma_ctrl_0_conduit_end.lcd_d_c_n
		lcd_dma_ctrl_0_conduit_end_lcd_wr_n    : out   std_logic;                                        --                                .lcd_wr_n
		lcd_dma_ctrl_0_conduit_end_lcd_data    : out   std_logic_vector(15 downto 0);                    --                                .lcd_data
		leds_external_connection_export_export : inout std_logic_vector(31 downto 0) := (others => '0'); -- leds_external_connection_export.export
		reset_reset_n                          : in    std_logic                     := '0';             --                           reset.reset_n
		sdram_controller_wire_addr             : out   std_logic_vector(11 downto 0);                    --           sdram_controller_wire.addr
		sdram_controller_wire_ba               : out   std_logic_vector(1 downto 0);                     --                                .ba
		sdram_controller_wire_cas_n            : out   std_logic;                                        --                                .cas_n
		sdram_controller_wire_cke              : out   std_logic;                                        --                                .cke
		sdram_controller_wire_cs_n             : out   std_logic;                                        --                                .cs_n
		sdram_controller_wire_dq               : inout std_logic_vector(15 downto 0) := (others => '0'); --                                .dq
		sdram_controller_wire_dqm              : out   std_logic_vector(1 downto 0);                     --                                .dqm
		sdram_controller_wire_ras_n            : out   std_logic;                                        --                                .ras_n
		sdram_controller_wire_we_n             : out   std_logic                                         --                                .we_n
	);
end entity model;

architecture rtl of model is
	component model_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(25 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component model_CPU;

	component DMA_LCD_ctrl is
		generic (
			SIZEOFINT16     : integer := 16;
			SIZEOFINT32     : integer := 32;
			SIZEOFAVALONADD : integer := 3
		);
		port (
			LCD_D_C_n_o              : out std_logic;                                        -- lcd_d_c_n
			LCD_WR_n_o               : out std_logic;                                        -- lcd_wr_n
			LCD_data_o               : out std_logic_vector(15 downto 0);                    -- lcd_data
			clk_i                    : in  std_logic                     := 'X';             -- clk
			reset_i                  : in  std_logic                     := 'X';             -- reset
			avalon_cs_i              : in  std_logic                     := 'X';             -- chipselect
			avalon_wr_i              : in  std_logic                     := 'X';             -- write
			avalon_rd_i              : in  std_logic                     := 'X';             -- read
			avalon_read_data_o       : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_address_i         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avalon_waitrequest_o     : out std_logic;                                        -- waitrequest
			avalon_write_data_i      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			master_address_o         : out std_logic_vector(31 downto 0);                    -- address
			master_read_o            : out std_logic;                                        -- read
			master_readdata_i        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			master_waitrequest_i     : in  std_logic                     := 'X';             -- waitrequest
			end_of_transaction_irq_o : out std_logic                                         -- irq
		);
	end component DMA_LCD_ctrl;

	component ParallelPort is
		port (
			Clk        : in    std_logic                     := 'X';             -- clk
			Address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			ChipSelect : in    std_logic                     := 'X';             -- chipselect
			Read       : in    std_logic                     := 'X';             -- read
			Write      : in    std_logic                     := 'X';             -- write
			ReadData   : out   std_logic_vector(31 downto 0);                    -- readdata
			WriteData  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nReset     : in    std_logic                     := 'X';             -- reset_n
			ParPort    : inout std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component ParallelPort;

	component model_SDRAM_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(22 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component model_SDRAM_controller;

	component model_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component model_jtag_uart;

	component model_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component model_sys_sdram_pll_0;

	component model_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component model_sysid_qsys_0;

	component model_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component model_timer_0;

	component model_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                           : in  std_logic                     := 'X';             -- clk
			LCD_DMA_CTRL_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                               : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                                  : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_readdatavalid                         : out std_logic;                                        -- readdatavalid
			CPU_data_master_write                                 : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address                        : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			LCD_DMA_CTRL_0_avalon_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			LCD_DMA_CTRL_0_avalon_master_waitrequest              : out std_logic;                                        -- waitrequest
			LCD_DMA_CTRL_0_avalon_master_read                     : in  std_logic                     := 'X';             -- read
			LCD_DMA_CTRL_0_avalon_master_readdata                 : out std_logic_vector(15 downto 0);                    -- readdata
			CPU_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                             : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                              : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			LCD_DMA_CTRL_0_avalon_slave_0_address                 : out std_logic_vector(2 downto 0);                     -- address
			LCD_DMA_CTRL_0_avalon_slave_0_write                   : out std_logic;                                        -- write
			LCD_DMA_CTRL_0_avalon_slave_0_read                    : out std_logic;                                        -- read
			LCD_DMA_CTRL_0_avalon_slave_0_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LCD_DMA_CTRL_0_avalon_slave_0_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			LCD_DMA_CTRL_0_avalon_slave_0_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			LCD_DMA_CTRL_0_avalon_slave_0_chipselect              : out std_logic;                                        -- chipselect
			LEDs_controller_0_avalon_slave_0_address              : out std_logic_vector(2 downto 0);                     -- address
			LEDs_controller_0_avalon_slave_0_write                : out std_logic;                                        -- write
			LEDs_controller_0_avalon_slave_0_read                 : out std_logic;                                        -- read
			LEDs_controller_0_avalon_slave_0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDs_controller_0_avalon_slave_0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			LEDs_controller_0_avalon_slave_0_chipselect           : out std_logic;                                        -- chipselect
			SDRAM_controller_s1_address                           : out std_logic_vector(22 downto 0);                    -- address
			SDRAM_controller_s1_write                             : out std_logic;                                        -- write
			SDRAM_controller_s1_read                              : out std_logic;                                        -- read
			SDRAM_controller_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_controller_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_controller_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_controller_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_controller_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_controller_s1_chipselect                        : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                    : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                      : out std_logic;                                        -- write
			timer_0_s1_readdata                                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                  : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                 : out std_logic                                         -- chipselect
		);
	end component model_mm_interconnect_0;

	component model_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component model_irq_mapper;

	component model_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component model_rst_controller;

	component model_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component model_rst_controller_001;

	signal sys_sdram_pll_0_sys_clk_clk                                   : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [CPU:clk, LCD_DMA_CTRL_0:clk_i, LEDs_controller_0:Clk, SDRAM_controller:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, rst_controller:clk, sysid_qsys_0:clock, timer_0:clk]
	signal lcd_dma_ctrl_0_avalon_master_readdata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_master_readdata -> LCD_DMA_CTRL_0:master_readdata_i
	signal lcd_dma_ctrl_0_avalon_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_master_waitrequest -> LCD_DMA_CTRL_0:master_waitrequest_i
	signal lcd_dma_ctrl_0_avalon_master_address                          : std_logic_vector(31 downto 0); -- LCD_DMA_CTRL_0:master_address_o -> mm_interconnect_0:LCD_DMA_CTRL_0_avalon_master_address
	signal lcd_dma_ctrl_0_avalon_master_read                             : std_logic;                     -- LCD_DMA_CTRL_0:master_read_o -> mm_interconnect_0:LCD_DMA_CTRL_0_avalon_master_read
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(25 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	signal cpu_data_master_write                                         : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(25 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_chipselect              : std_logic;                     -- mm_interconnect_0:SDRAM_controller_s1_chipselect -> SDRAM_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                : std_logic_vector(15 downto 0); -- SDRAM_controller:za_data -> mm_interconnect_0:SDRAM_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest             : std_logic;                     -- SDRAM_controller:za_waitrequest -> mm_interconnect_0:SDRAM_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                 : std_logic_vector(22 downto 0); -- mm_interconnect_0:SDRAM_controller_s1_address -> SDRAM_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                    : std_logic;                     -- mm_interconnect_0:SDRAM_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid           : std_logic;                     -- SDRAM_controller:za_valid -> mm_interconnect_0:SDRAM_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                   : std_logic;                     -- mm_interconnect_0:SDRAM_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata               : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_controller_s1_writedata -> SDRAM_controller:az_data
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:LEDs_controller_0_avalon_slave_0_chipselect -> LEDs_controller_0:ChipSelect
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_readdata   : std_logic_vector(31 downto 0); -- LEDs_controller_0:ReadData -> mm_interconnect_0:LEDs_controller_0_avalon_slave_0_readdata
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_address    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:LEDs_controller_0_avalon_slave_0_address -> LEDs_controller_0:Address
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:LEDs_controller_0_avalon_slave_0_read -> LEDs_controller_0:Read
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:LEDs_controller_0_avalon_slave_0_write -> LEDs_controller_0:Write
	signal mm_interconnect_0_leds_controller_0_avalon_slave_0_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDs_controller_0_avalon_slave_0_writedata -> LEDs_controller_0:WriteData
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_chipselect    : std_logic;                     -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_chipselect -> LCD_DMA_CTRL_0:avalon_cs_i
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_readdata      : std_logic_vector(31 downto 0); -- LCD_DMA_CTRL_0:avalon_read_data_o -> mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_readdata
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_waitrequest   : std_logic;                     -- LCD_DMA_CTRL_0:avalon_waitrequest_o -> mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_address       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_address -> LCD_DMA_CTRL_0:avalon_address_i
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_read          : std_logic;                     -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_read -> LCD_DMA_CTRL_0:avalon_rd_i
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_write         : std_logic;                     -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_write -> LCD_DMA_CTRL_0:avalon_wr_i
	signal mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_DMA_CTRL_0_avalon_slave_0_writedata -> LCD_DMA_CTRL_0:avalon_write_data_i
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata         : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_timer_0_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                         : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                            : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- LCD_DMA_CTRL_0:end_of_transaction_irq_o -> irq_mapper:receiver2_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [LCD_DMA_CTRL_0:reset_i, irq_mapper:reset, mm_interconnect_0:LCD_DMA_CTRL_0_reset_sink_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                 : std_logic;                     -- CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> sys_sdram_pll_0:ref_reset_reset
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv          : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> SDRAM_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> SDRAM_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> SDRAM_controller:az_wr_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, LEDs_controller_0:nReset, SDRAM_controller:reset_n, jtag_uart:rst_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	cpu : component model_CPU
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                       --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	lcd_dma_ctrl_0 : component DMA_LCD_ctrl
		generic map (
			SIZEOFINT16     => 16,
			SIZEOFINT32     => 32,
			SIZEOFAVALONADD => 3
		)
		port map (
			LCD_D_C_n_o              => lcd_dma_ctrl_0_conduit_end_lcd_d_c_n,                        --    conduit_end.lcd_d_c_n
			LCD_WR_n_o               => lcd_dma_ctrl_0_conduit_end_lcd_wr_n,                         --               .lcd_wr_n
			LCD_data_o               => lcd_dma_ctrl_0_conduit_end_lcd_data,                         --               .lcd_data
			clk_i                    => sys_sdram_pll_0_sys_clk_clk,                                 --     clock_sink.clk
			reset_i                  => rst_controller_reset_out_reset,                              --     reset_sink.reset
			avalon_cs_i              => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_chipselect,  -- avalon_slave_0.chipselect
			avalon_wr_i              => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_write,       --               .write
			avalon_rd_i              => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_read,        --               .read
			avalon_read_data_o       => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_readdata,    --               .readdata
			avalon_address_i         => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_address,     --               .address
			avalon_waitrequest_o     => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_waitrequest, --               .waitrequest
			avalon_write_data_i      => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_writedata,   --               .writedata
			master_address_o         => lcd_dma_ctrl_0_avalon_master_address,                        --  avalon_master.address
			master_read_o            => lcd_dma_ctrl_0_avalon_master_read,                           --               .read
			master_readdata_i        => lcd_dma_ctrl_0_avalon_master_readdata,                       --               .readdata
			master_waitrequest_i     => lcd_dma_ctrl_0_avalon_master_waitrequest,                    --               .waitrequest
			end_of_transaction_irq_o => irq_mapper_receiver2_irq                                     --            irq.irq
		);

	leds_controller_0 : component ParallelPort
		port map (
			Clk        => sys_sdram_pll_0_sys_clk_clk,                                   --          clock.clk
			Address    => mm_interconnect_0_leds_controller_0_avalon_slave_0_address,    -- avalon_slave_0.address
			ChipSelect => mm_interconnect_0_leds_controller_0_avalon_slave_0_chipselect, --               .chipselect
			Read       => mm_interconnect_0_leds_controller_0_avalon_slave_0_read,       --               .read
			Write      => mm_interconnect_0_leds_controller_0_avalon_slave_0_write,      --               .write
			ReadData   => mm_interconnect_0_leds_controller_0_avalon_slave_0_readdata,   --               .readdata
			WriteData  => mm_interconnect_0_leds_controller_0_avalon_slave_0_writedata,  --               .writedata
			nReset     => rst_controller_reset_out_reset_ports_inv,                      --     reset_sink.reset_n
			ParPort    => leds_external_connection_export_export                         --  conduit_end_1.export
		);

	sdram_controller : component model_SDRAM_controller
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_wire_we_n                                  --      .export
		);

	jtag_uart : component model_jtag_uart
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	sys_sdram_pll_0 : component model_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			reset_source_reset => open                                -- reset_source.reset
		);

	sysid_qsys_0 : component model_sysid_qsys_0
		port map (
			clock    => sys_sdram_pll_0_sys_clk_clk,                             --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component model_timer_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component model_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                           => sys_sdram_pll_0_sys_clk_clk,                                   --                         sys_sdram_pll_0_sys_clk.clk
			LCD_DMA_CTRL_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                -- LCD_DMA_CTRL_0_reset_sink_reset_bridge_in_reset.reset
			CPU_data_master_address                               => cpu_data_master_address,                                       --                                 CPU_data_master.address
			CPU_data_master_waitrequest                           => cpu_data_master_waitrequest,                                   --                                                .waitrequest
			CPU_data_master_byteenable                            => cpu_data_master_byteenable,                                    --                                                .byteenable
			CPU_data_master_read                                  => cpu_data_master_read,                                          --                                                .read
			CPU_data_master_readdata                              => cpu_data_master_readdata,                                      --                                                .readdata
			CPU_data_master_readdatavalid                         => cpu_data_master_readdatavalid,                                 --                                                .readdatavalid
			CPU_data_master_write                                 => cpu_data_master_write,                                         --                                                .write
			CPU_data_master_writedata                             => cpu_data_master_writedata,                                     --                                                .writedata
			CPU_data_master_debugaccess                           => cpu_data_master_debugaccess,                                   --                                                .debugaccess
			CPU_instruction_master_address                        => cpu_instruction_master_address,                                --                          CPU_instruction_master.address
			CPU_instruction_master_waitrequest                    => cpu_instruction_master_waitrequest,                            --                                                .waitrequest
			CPU_instruction_master_read                           => cpu_instruction_master_read,                                   --                                                .read
			CPU_instruction_master_readdata                       => cpu_instruction_master_readdata,                               --                                                .readdata
			CPU_instruction_master_readdatavalid                  => cpu_instruction_master_readdatavalid,                          --                                                .readdatavalid
			LCD_DMA_CTRL_0_avalon_master_address                  => lcd_dma_ctrl_0_avalon_master_address,                          --                    LCD_DMA_CTRL_0_avalon_master.address
			LCD_DMA_CTRL_0_avalon_master_waitrequest              => lcd_dma_ctrl_0_avalon_master_waitrequest,                      --                                                .waitrequest
			LCD_DMA_CTRL_0_avalon_master_read                     => lcd_dma_ctrl_0_avalon_master_read,                             --                                                .read
			LCD_DMA_CTRL_0_avalon_master_readdata                 => lcd_dma_ctrl_0_avalon_master_readdata,                         --                                                .readdata
			CPU_debug_mem_slave_address                           => mm_interconnect_0_cpu_debug_mem_slave_address,                 --                             CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                             => mm_interconnect_0_cpu_debug_mem_slave_write,                   --                                                .write
			CPU_debug_mem_slave_read                              => mm_interconnect_0_cpu_debug_mem_slave_read,                    --                                                .read
			CPU_debug_mem_slave_readdata                          => mm_interconnect_0_cpu_debug_mem_slave_readdata,                --                                                .readdata
			CPU_debug_mem_slave_writedata                         => mm_interconnect_0_cpu_debug_mem_slave_writedata,               --                                                .writedata
			CPU_debug_mem_slave_byteenable                        => mm_interconnect_0_cpu_debug_mem_slave_byteenable,              --                                                .byteenable
			CPU_debug_mem_slave_waitrequest                       => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,             --                                                .waitrequest
			CPU_debug_mem_slave_debugaccess                       => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,             --                                                .debugaccess
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,         --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,           --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,            --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      --                                                .chipselect
			LCD_DMA_CTRL_0_avalon_slave_0_address                 => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_address,       --                   LCD_DMA_CTRL_0_avalon_slave_0.address
			LCD_DMA_CTRL_0_avalon_slave_0_write                   => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_write,         --                                                .write
			LCD_DMA_CTRL_0_avalon_slave_0_read                    => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_read,          --                                                .read
			LCD_DMA_CTRL_0_avalon_slave_0_readdata                => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_readdata,      --                                                .readdata
			LCD_DMA_CTRL_0_avalon_slave_0_writedata               => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_writedata,     --                                                .writedata
			LCD_DMA_CTRL_0_avalon_slave_0_waitrequest             => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_waitrequest,   --                                                .waitrequest
			LCD_DMA_CTRL_0_avalon_slave_0_chipselect              => mm_interconnect_0_lcd_dma_ctrl_0_avalon_slave_0_chipselect,    --                                                .chipselect
			LEDs_controller_0_avalon_slave_0_address              => mm_interconnect_0_leds_controller_0_avalon_slave_0_address,    --                LEDs_controller_0_avalon_slave_0.address
			LEDs_controller_0_avalon_slave_0_write                => mm_interconnect_0_leds_controller_0_avalon_slave_0_write,      --                                                .write
			LEDs_controller_0_avalon_slave_0_read                 => mm_interconnect_0_leds_controller_0_avalon_slave_0_read,       --                                                .read
			LEDs_controller_0_avalon_slave_0_readdata             => mm_interconnect_0_leds_controller_0_avalon_slave_0_readdata,   --                                                .readdata
			LEDs_controller_0_avalon_slave_0_writedata            => mm_interconnect_0_leds_controller_0_avalon_slave_0_writedata,  --                                                .writedata
			LEDs_controller_0_avalon_slave_0_chipselect           => mm_interconnect_0_leds_controller_0_avalon_slave_0_chipselect, --                                                .chipselect
			SDRAM_controller_s1_address                           => mm_interconnect_0_sdram_controller_s1_address,                 --                             SDRAM_controller_s1.address
			SDRAM_controller_s1_write                             => mm_interconnect_0_sdram_controller_s1_write,                   --                                                .write
			SDRAM_controller_s1_read                              => mm_interconnect_0_sdram_controller_s1_read,                    --                                                .read
			SDRAM_controller_s1_readdata                          => mm_interconnect_0_sdram_controller_s1_readdata,                --                                                .readdata
			SDRAM_controller_s1_writedata                         => mm_interconnect_0_sdram_controller_s1_writedata,               --                                                .writedata
			SDRAM_controller_s1_byteenable                        => mm_interconnect_0_sdram_controller_s1_byteenable,              --                                                .byteenable
			SDRAM_controller_s1_readdatavalid                     => mm_interconnect_0_sdram_controller_s1_readdatavalid,           --                                                .readdatavalid
			SDRAM_controller_s1_waitrequest                       => mm_interconnect_0_sdram_controller_s1_waitrequest,             --                                                .waitrequest
			SDRAM_controller_s1_chipselect                        => mm_interconnect_0_sdram_controller_s1_chipselect,              --                                                .chipselect
			sysid_qsys_0_control_slave_address                    => mm_interconnect_0_sysid_qsys_0_control_slave_address,          --                      sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                   => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,         --                                                .readdata
			timer_0_s1_address                                    => mm_interconnect_0_timer_0_s1_address,                          --                                      timer_0_s1.address
			timer_0_s1_write                                      => mm_interconnect_0_timer_0_s1_write,                            --                                                .write
			timer_0_s1_readdata                                   => mm_interconnect_0_timer_0_s1_readdata,                         --                                                .readdata
			timer_0_s1_writedata                                  => mm_interconnect_0_timer_0_s1_writedata,                        --                                                .writedata
			timer_0_s1_chipselect                                 => mm_interconnect_0_timer_0_s1_chipselect                        --                                                .chipselect
		);

	irq_mapper : component model_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component model_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component model_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of model
